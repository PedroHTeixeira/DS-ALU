----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:	14:44:37 05/19/2022
-- Design Name:
-- Module Name:	ADDER - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ADDER is
	Port ( x : in  STD_LOGIC;
       	y : in  STD_LOGIC;
       	cin : in  STD_LOGIC;
       	cout : out  STD_LOGIC;
       	z : out  STD_LOGIC);
end ADDER;

architecture Behavioral of ADDER is

begin
    z <= (x XOR y) XOR cin;
    cout <= (x AND y) OR (cin AND (x XOR y));

end Behavioral;
